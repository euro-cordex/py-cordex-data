netcdf tas_EUR-11_ECMWF-ERAINT_evaluation_r1i1p1_GERICS-REMO2015_v1_mon_198001-198012 {
dimensions:
	time = UNLIMITED ; // (12 currently)
	bnds = 2 ;
	rlon = 424 ;
	rlat = 412 ;
	vertices = 4 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1949-12-01T00:00:00Z" ;
		time:calendar = "proleptic_gregorian" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;
	float lon(rlat, rlon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude coordinate" ;
		lon:units = "degrees_east" ;
		lon:_CoordinateAxisType = "Lon" ;
		lon:bounds = "lon_bnds" ;
	float lon_bnds(rlat, rlon, vertices) ;
	float lat(rlat, rlon) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude coordinate" ;
		lat:units = "degrees_north" ;
		lat:_CoordinateAxisType = "Lat" ;
		lat:bounds = "lat_bnds" ;
	float lat_bnds(rlat, rlon, vertices) ;
	double rlon(rlon) ;
		rlon:standard_name = "grid_longitude" ;
		rlon:long_name = "longitude in rotated pole grid" ;
		rlon:units = "degrees" ;
		rlon:axis = "X" ;
	double rlat(rlat) ;
		rlat:standard_name = "grid_latitude" ;
		rlat:long_name = "latitude in rotated pole grid" ;
		rlat:units = "degrees" ;
		rlat:axis = "Y" ;
	int rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:grid_north_pole_latitude = 39.25 ;
		rotated_latitude_longitude:grid_north_pole_longitude = -162. ;
		rotated_latitude_longitude:north_pole_grid_longitude = 0. ;
	double height ;
		height:standard_name = "height" ;
		height:long_name = "height" ;
		height:units = "m" ;
		height:positive = "up" ;
		height:axis = "Z" ;
	float tas(time, rlat, rlon) ;
		tas:standard_name = "air_temperature" ;
		tas:long_name = "Near-Surface Air Temperature" ;
		tas:units = "K" ;
		tas:grid_mapping = "rotated_latitude_longitude" ;
		tas:coordinates = "height lat lon" ;
		tas:_FillValue = 1.e+20f ;
		tas:missing_value = 1.e+20f ;
		tas:comment = "daily-mean near-surface (usually, 2 meter) air temperature." ;
		tas:cell_methods = "time: mean" ;
		tas:history = "2018-06-15T15:20:54Z altered by CMOR: Treated scalar dimension: \'height\'." ;
		tas:associated_files = "gridspecFile: gridspec_atmos_fx_GERICS-REMO2015_evaluation_r0i0p0.nc" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.6.1|hdf5libversion=1.8.14" ;
		:CDI = "Climate Data Interface version 1.9.7.1 (http://mpimet.mpg.de/cdi)" ;
		:history = "Thu Nov 25 12:23:50 2021: cdo selyear,1980 tas_EUR-11_ECMWF-ERAINT_evaluation_r1i1p1_GERICS-REMO2015_v1_mon_197902-198012.nc tas_EUR-11_ECMWF-ERAINT_evaluation_r1i1p1_GERICS-REMO2015_v1_mon_198001-198012.nc\n",
			"2018-06-15T15:20:54Z CMOR rewrote data to comply with CF standards and CORDEX requirements." ;
		:source = "GERICS-REMO2015" ;
		:institution = "Helmholtz-Zentrum Geesthacht, Climate Service Center Germany" ;
		:Conventions = "CF-1.4" ;
		:institute_id = "GERICS" ;
		:experiment_id = "evaluation" ;
		:model_id = "GERICS-REMO2015" ;
		:contact = "gerics-cordex@hzg.de" ;
		:comment = "CORDEX Europe RCM REMO 0.11 deg EUR-11." ;
		:references = "http://www.remo-rcm.de/" ;
		:initialization_method = 1 ;
		:physics_version = 1 ;
		:tracking_id = "07c8a6b9-424a-4867-815c-5fbce2675d0b" ;
		:CORDEX_domain = "EUR-11" ;
		:driving_experiment = "ECMWF-ERAINT, evaluation, r1i1p1" ;
		:driving_model_id = "ECMWF-ERAINT" ;
		:driving_model_ensemble_member = "r1i1p1" ;
		:driving_experiment_name = "evaluation" ;
		:rcm_version_id = "v1" ;
		:product = "output" ;
		:experiment = "Evaluation run with reanalysis forcing" ;
		:frequency = "mon" ;
		:creation_date = "2018-06-15T15:20:54Z" ;
		:project_id = "CORDEX" ;
		:table_id = "Table mon (Mar 2015) db0b230ff4a2c922671f0c21978b6242" ;
		:title = "GERICS-REMO2015 model output prepared for CORDEX Evaluation run with reanalysis forcing" ;
		:modeling_realm = "atmos" ;
		:realization = 1 ;
		:cmor_version = "2.9.1" ;
		:CDO = "Climate Data Operators version 1.9.7.1 (http://mpimet.mpg.de/cdo)" ;
data:

 time = 11003.5, 11033.5, 11063.5, 11094, 11124.5, 11155, 11185.5, 11216.5, 
    11247, 11277.5, 11308, 11338.5 ;

 time_bnds =
  10988, 11019,
  11019, 11048,
  11048, 11079,
  11079, 11109,
  11109, 11140,
  11140, 11170,
  11170, 11201,
  11201, 11232,
  11232, 11262,
  11262, 11293,
  11293, 11323,
  11323, 11354 ;

 rlon = -28.375, -28.265, -28.155, -28.045, -27.935, -27.825, -27.715, 
    -27.605, -27.495, -27.385, -27.275, -27.165, -27.055, -26.945, -26.835, 
    -26.725, -26.615, -26.505, -26.395, -26.285, -26.175, -26.065, -25.955, 
    -25.845, -25.735, -25.625, -25.515, -25.405, -25.295, -25.185, -25.075, 
    -24.965, -24.855, -24.745, -24.635, -24.525, -24.415, -24.305, -24.195, 
    -24.085, -23.975, -23.865, -23.755, -23.645, -23.535, -23.425, -23.315, 
    -23.205, -23.095, -22.985, -22.875, -22.765, -22.655, -22.545, -22.435, 
    -22.325, -22.215, -22.105, -21.995, -21.885, -21.775, -21.665, -21.555, 
    -21.445, -21.335, -21.225, -21.115, -21.005, -20.895, -20.785, -20.675, 
    -20.565, -20.455, -20.345, -20.235, -20.125, -20.015, -19.905, -19.795, 
    -19.685, -19.575, -19.465, -19.355, -19.245, -19.135, -19.025, -18.915, 
    -18.805, -18.695, -18.585, -18.475, -18.365, -18.255, -18.145, -18.035, 
    -17.925, -17.815, -17.705, -17.595, -17.485, -17.375, -17.265, -17.155, 
    -17.045, -16.935, -16.825, -16.715, -16.605, -16.495, -16.385, -16.275, 
    -16.165, -16.055, -15.945, -15.835, -15.725, -15.615, -15.505, -15.395, 
    -15.285, -15.175, -15.065, -14.955, -14.845, -14.735, -14.625, -14.515, 
    -14.405, -14.295, -14.185, -14.075, -13.965, -13.855, -13.745, -13.635, 
    -13.525, -13.415, -13.305, -13.195, -13.085, -12.975, -12.865, -12.755, 
    -12.645, -12.535, -12.425, -12.315, -12.205, -12.095, -11.985, -11.875, 
    -11.765, -11.655, -11.545, -11.435, -11.325, -11.215, -11.105, -10.995, 
    -10.885, -10.775, -10.665, -10.555, -10.445, -10.335, -10.225, -10.115, 
    -10.005, -9.895, -9.785, -9.675, -9.565, -9.455, -9.345, -9.235, -9.125, 
    -9.015, -8.905, -8.795, -8.685, -8.575, -8.465, -8.355, -8.245, -8.135, 
    -8.025, -7.915, -7.805, -7.695, -7.585, -7.475, -7.365, -7.255, -7.145, 
    -7.035, -6.925, -6.815, -6.705, -6.595, -6.485, -6.375, -6.265, -6.155, 
    -6.045, -5.935, -5.825, -5.715, -5.605, -5.495, -5.385, -5.275, -5.165, 
    -5.055, -4.945, -4.835, -4.725, -4.615, -4.505, -4.395, -4.285, -4.175, 
    -4.065, -3.955, -3.845, -3.735, -3.625, -3.515, -3.405, -3.295, -3.185, 
    -3.075, -2.965, -2.855, -2.745, -2.635, -2.525, -2.415, -2.305, -2.195, 
    -2.085, -1.975, -1.865, -1.755, -1.645, -1.535, -1.425, -1.315, -1.205, 
    -1.095, -0.985000000000001, -0.875000000000001, -0.765000000000001, 
    -0.655000000000001, -0.545000000000001, -0.435000000000001, 
    -0.325000000000001, -0.215000000000001, -0.105000000000001, 
    0.00499999999999944, 0.114999999999999, 0.224999999999999, 
    0.334999999999999, 0.444999999999999, 0.554999999999999, 
    0.664999999999999, 0.774999999999999, 0.884999999999999, 
    0.994999999999999, 1.105, 1.215, 1.325, 1.435, 1.545, 1.655, 1.765, 
    1.875, 1.985, 2.095, 2.205, 2.315, 2.425, 2.535, 2.645, 2.755, 2.865, 
    2.975, 3.085, 3.195, 3.305, 3.415, 3.525, 3.635, 3.745, 3.855, 3.965, 
    4.075, 4.185, 4.295, 4.405, 4.515, 4.625, 4.735, 4.845, 4.955, 5.065, 
    5.175, 5.285, 5.395, 5.505, 5.615, 5.725, 5.835, 5.945, 6.055, 6.165, 
    6.275, 6.385, 6.495, 6.605, 6.715, 6.825, 6.935, 7.045, 7.155, 7.265, 
    7.375, 7.485, 7.595, 7.705, 7.815, 7.925, 8.035, 8.145, 8.255, 8.365, 
    8.475, 8.585, 8.695, 8.805, 8.915, 9.025, 9.135, 9.245, 9.355, 9.465, 
    9.575, 9.685, 9.795, 9.905, 10.015, 10.125, 10.235, 10.345, 10.455, 
    10.565, 10.675, 10.785, 10.895, 11.005, 11.115, 11.225, 11.335, 11.445, 
    11.555, 11.665, 11.775, 11.885, 11.995, 12.105, 12.215, 12.325, 12.435, 
    12.545, 12.655, 12.765, 12.875, 12.985, 13.095, 13.205, 13.315, 13.425, 
    13.535, 13.645, 13.755, 13.865, 13.975, 14.085, 14.195, 14.305, 14.415, 
    14.525, 14.635, 14.745, 14.855, 14.965, 15.075, 15.185, 15.295, 15.405, 
    15.515, 15.625, 15.735, 15.845, 15.955, 16.065, 16.175, 16.285, 16.395, 
    16.505, 16.615, 16.725, 16.835, 16.945, 17.055, 17.165, 17.275, 17.385, 
    17.495, 17.605, 17.715, 17.825, 17.935, 18.045, 18.155 ;

 rlat = -23.375, -23.265, -23.155, -23.045, -22.935, -22.825, -22.715, 
    -22.605, -22.495, -22.385, -22.275, -22.165, -22.055, -21.945, -21.835, 
    -21.725, -21.615, -21.505, -21.395, -21.285, -21.175, -21.065, -20.955, 
    -20.845, -20.735, -20.625, -20.515, -20.405, -20.295, -20.185, -20.075, 
    -19.965, -19.855, -19.745, -19.635, -19.525, -19.415, -19.305, -19.195, 
    -19.085, -18.975, -18.865, -18.755, -18.645, -18.535, -18.425, -18.315, 
    -18.205, -18.095, -17.985, -17.875, -17.765, -17.655, -17.545, -17.435, 
    -17.325, -17.215, -17.105, -16.995, -16.885, -16.775, -16.665, -16.555, 
    -16.445, -16.335, -16.225, -16.115, -16.005, -15.895, -15.785, -15.675, 
    -15.565, -15.455, -15.345, -15.235, -15.125, -15.015, -14.905, -14.795, 
    -14.685, -14.575, -14.465, -14.355, -14.245, -14.135, -14.025, -13.915, 
    -13.805, -13.695, -13.585, -13.475, -13.365, -13.255, -13.145, -13.035, 
    -12.925, -12.815, -12.705, -12.595, -12.485, -12.375, -12.265, -12.155, 
    -12.045, -11.935, -11.825, -11.715, -11.605, -11.495, -11.385, -11.275, 
    -11.165, -11.055, -10.945, -10.835, -10.725, -10.615, -10.505, -10.395, 
    -10.285, -10.175, -10.065, -9.955, -9.845, -9.735, -9.625, -9.515, 
    -9.405, -9.295, -9.185, -9.075, -8.965, -8.855, -8.745, -8.635, -8.525, 
    -8.415, -8.305, -8.195, -8.085, -7.975, -7.865, -7.755, -7.645, -7.535, 
    -7.425, -7.315, -7.205, -7.095, -6.985, -6.875, -6.765, -6.655, -6.545, 
    -6.435, -6.325, -6.215, -6.105, -5.995, -5.885, -5.775, -5.665, -5.555, 
    -5.445, -5.335, -5.225, -5.115, -5.005, -4.895, -4.785, -4.675, -4.565, 
    -4.455, -4.345, -4.235, -4.125, -4.015, -3.905, -3.795, -3.685, -3.575, 
    -3.465, -3.355, -3.245, -3.135, -3.025, -2.915, -2.805, -2.695, -2.585, 
    -2.475, -2.365, -2.255, -2.145, -2.035, -1.925, -1.815, -1.705, -1.595, 
    -1.485, -1.375, -1.265, -1.155, -1.045, -0.935000000000001, 
    -0.825000000000001, -0.715000000000001, -0.605000000000001, 
    -0.495000000000001, -0.385000000000001, -0.275000000000001, 
    -0.165000000000001, -0.0550000000000006, 0.0549999999999994, 
    0.164999999999999, 0.274999999999999, 0.384999999999999, 
    0.494999999999999, 0.604999999999999, 0.714999999999999, 
    0.824999999999999, 0.934999999999999, 1.045, 1.155, 1.265, 1.375, 1.485, 
    1.595, 1.705, 1.815, 1.925, 2.035, 2.145, 2.255, 2.365, 2.475, 2.585, 
    2.695, 2.805, 2.915, 3.025, 3.135, 3.245, 3.355, 3.465, 3.575, 3.685, 
    3.795, 3.905, 4.015, 4.125, 4.235, 4.345, 4.455, 4.565, 4.675, 4.785, 
    4.895, 5.005, 5.115, 5.225, 5.335, 5.445, 5.555, 5.665, 5.775, 5.885, 
    5.995, 6.105, 6.215, 6.325, 6.435, 6.545, 6.655, 6.765, 6.875, 6.985, 
    7.095, 7.205, 7.315, 7.425, 7.535, 7.645, 7.755, 7.865, 7.975, 8.085, 
    8.195, 8.305, 8.415, 8.525, 8.635, 8.745, 8.855, 8.965, 9.075, 9.185, 
    9.295, 9.405, 9.515, 9.625, 9.735, 9.845, 9.955, 10.065, 10.175, 10.285, 
    10.395, 10.505, 10.615, 10.725, 10.835, 10.945, 11.055, 11.165, 11.275, 
    11.385, 11.495, 11.605, 11.715, 11.825, 11.935, 12.045, 12.155, 12.265, 
    12.375, 12.485, 12.595, 12.705, 12.815, 12.925, 13.035, 13.145, 13.255, 
    13.365, 13.475, 13.585, 13.695, 13.805, 13.915, 14.025, 14.135, 14.245, 
    14.355, 14.465, 14.575, 14.685, 14.795, 14.905, 15.015, 15.125, 15.235, 
    15.345, 15.455, 15.565, 15.675, 15.785, 15.895, 16.005, 16.115, 16.225, 
    16.335, 16.445, 16.555, 16.665, 16.775, 16.885, 16.995, 17.105, 17.215, 
    17.325, 17.435, 17.545, 17.655, 17.765, 17.875, 17.985, 18.095, 18.205, 
    18.315, 18.425, 18.535, 18.645, 18.755, 18.865, 18.975, 19.085, 19.195, 
    19.305, 19.415, 19.525, 19.635, 19.745, 19.855, 19.965, 20.075, 20.185, 
    20.295, 20.405, 20.515, 20.625, 20.735, 20.845, 20.955, 21.065, 21.175, 
    21.285, 21.395, 21.505, 21.615, 21.725, 21.835 ;
}
